/**
* This module implements a decoder for handling the requests given to the FPGA. The handling is
* based on the established communication protocol found in - (LINK).
*/
module RequestHandler ();

endmodule
