/**
* This module implements a high level facade for handling responses off up to 32 different sensors.
*
* NOTE: Currently only working with the DHT11 sensor, whose module is found in this project by the
* name of `DHT11.v`.
*/
module SensorDecoder ();

endmodule
